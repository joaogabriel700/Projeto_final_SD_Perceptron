library verilog;
use verilog.vl_types.all;
entity decoder_7seg_vlg_check_tst is
    port(
        s0              : in     vl_logic;
        s1              : in     vl_logic;
        s2              : in     vl_logic;
        s3              : in     vl_logic;
        s4              : in     vl_logic;
        s5              : in     vl_logic;
        s6              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decoder_7seg_vlg_check_tst;
