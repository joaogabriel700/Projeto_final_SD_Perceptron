library verilog;
use verilog.vl_types.all;
entity register_36_vlg_vec_tst is
end register_36_vlg_vec_tst;
