library verilog;
use verilog.vl_types.all;
entity multiplicador_completo_vlg_vec_tst is
end multiplicador_completo_vlg_vec_tst;
