library verilog;
use verilog.vl_types.all;
entity perceptron_vlg_vec_tst is
end perceptron_vlg_vec_tst;
