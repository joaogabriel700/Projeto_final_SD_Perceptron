entity multiplicador_completo is 
    port(
        in_a : in bit_vector(15 downto 0);
        in_b : in bit_vector(7 downto 0);
        resultado : out bit_vector(23 downto 0) 
    );
    end multiplicador_completo;

architecture behav of multiplicador_completo is 

component multiplicador_24bit is
    port(
        dados : in bit_vector(15 downto 0);
        inp : in bit_vector(7 downto 0);
        P: out bit_vector(23 downto 0)
    );
end component; 

component corretor_sinal is 
    port(
        entrada : in bit_vector(23 downto 0);
        comp : in bit;
        saida : out bit_vector( 23 downto 0)
    );
end component; 

signal sinal_a, sinal_b,sinal_f : bit;

signal A_ex : bit_vector(23 downto 0);
signal A_p  : bit_vector(23 downto 0);

signal B_ex : bit_vector(23 downto 0);
signal B_p : bit_vector(23 downto 0);

signal P_sem_sinal : bit_vector(23 downto 0); 

begin 

sinal_a <= in_a(15);

sinal_b <= in_b(7);

sinal_f <= sinal_a xor sinal_b; 

A_ex(15 downto 0) <= in_a;

A_ex(16) <=in_a(15);

A_ex(17) <=in_a(15);

A_ex(18) <=in_a(15);

A_ex(19) <=in_a(15);

A_ex(20) <=in_a(15);

A_ex(21) <=in_a(15);

A_ex(22) <=in_a(15);

A_ex(23) <=in_a(15);

B_ex(7 downto 0) <= in_b;

B_ex(8) <= in_b(7);

B_ex(9) <= in_b(7); 

B_ex(10) <= in_b(7); 

B_ex(11) <= in_b(7); 

B_ex(12) <= in_b(7); 

B_ex(13) <= in_b(7); 

B_ex(14) <= in_b(7); 

B_ex(15) <= in_b(7); 

B_ex(16) <= in_b(7); 

B_ex(17) <= in_b(7); 

B_ex(18) <= in_b(7); 

B_ex(19) <= in_b(7);

B_ex(20) <= in_b(7); 

B_ex(21) <= in_b(7); 

B_ex(22) <= in_b(7); 

B_ex(23) <= in_b(7); 

corrige_a: corretor_sinal port map(
            entrada => A_ex,
            comp => sinal_a,
            saida => A_p
);

corrige_b : corretor_sinal port map(
            entrada => B_ex,
            comp => sinal_b,
            saida => B_p
);

multiplica : multiplicador_24bit port map(
            dados => A_p(15 downto 0),
            inp => B_p(7 downto 0),
            P => P_sem_sinal
);

corrige_saida : corretor_sinal port map(
            entrada => P_sem_sinal,
            comp => sinal_f,
            saida => resultado
);

end architecture behav;