library verilog;
use verilog.vl_types.all;
entity decoder_7seg_vlg_sample_tst is
    port(
        into            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end decoder_7seg_vlg_sample_tst;
