library verilog;
use verilog.vl_types.all;
entity mux_4x1_24bit_vlg_vec_tst is
end mux_4x1_24bit_vlg_vec_tst;
