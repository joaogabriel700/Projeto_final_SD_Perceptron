library verilog;
use verilog.vl_types.all;
entity rom_3x16_vlg_vec_tst is
end rom_3x16_vlg_vec_tst;
