library verilog;
use verilog.vl_types.all;
entity somador_24bit_vlg_check_tst is
    port(
        S               : in     vl_logic_vector(23 downto 0);
        sampler_rx      : in     vl_logic
    );
end somador_24bit_vlg_check_tst;
