library verilog;
use verilog.vl_types.all;
entity multiplicador_24bit_vlg_vec_tst is
end multiplicador_24bit_vlg_vec_tst;
