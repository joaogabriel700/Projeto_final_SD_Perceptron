library verilog;
use verilog.vl_types.all;
entity somador_24bit_vlg_vec_tst is
end somador_24bit_vlg_vec_tst;
