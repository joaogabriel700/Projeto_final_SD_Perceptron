library verilog;
use verilog.vl_types.all;
entity multiplicador_24bit_vlg_check_tst is
    port(
        P               : in     vl_logic_vector(23 downto 0);
        sampler_rx      : in     vl_logic
    );
end multiplicador_24bit_vlg_check_tst;
